`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/06/2022 05:26:28 PM
// Design Name: 
// Module Name: binary_to_number
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bcd_to_number(
    input [3:0] hours0,hours1, minutes0,minutes1, seconds0,seconds1, milliseconds0,milliseconds1,milliseconds2,
    output reg [13:0] h, m, s,
    output reg [20:0] k
    );
    always@(*)begin
        case (hours1)
            4'b0000: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1111101;
            4'b0001: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1100000;
            4'b0010: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b0110111;
            4'b0011: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1100111;
            4'b0100: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1101010;
            4'b0101: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1001111;
            4'b0110: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1011111;
            4'b0111: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1100001;
            4'b1000: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1111111;
            4'b1001: {h[6],h[5],h[4],h[3],h[2],h[1],h[0]}=7'b1101011;
        endcase
        case(hours0)
            4'b0000: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1111101;
            4'b0001: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1100000;
            4'b0010: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b0110111;
            4'b0011: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1100111;
            4'b0100: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1101010;
            4'b0101: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1001111;
            4'b0110: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1011111;
            4'b0111: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1100001;
            4'b1000: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1111111;
            4'b1001: {h[13],h[12],h[11],h[10],h[9],h[8],h[7]}=7'b1101011; 
        endcase
        case(minutes1)
            4'b0000: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1111101;
            4'b0001: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1100000; 
            4'b0010: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b0110111;
            4'b0011: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1100111;
            4'b0100: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1101010;
            4'b0101: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1001111;
            /*
            4'b0110: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1111100;
            4'b0111: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1000011;
            4'b1000: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1111111;
            4'b1001: {m[6],m[5],m[4],m[3],m[2],m[1],m[0]}=7'b1101011; 
            */
        endcase
        case(minutes0)
            4'b0000: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1111101;
            4'b0001: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1100000; 
            4'b0010: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b0110111;
            4'b0011: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1100111;
            4'b0100: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1101010;
            4'b0101: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1001111;
            4'b0110: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1011111;
            4'b0111: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1100001;
            4'b1000: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1111111;
            4'b1001: {m[13],m[12],m[11],m[10],m[9],m[8],m[7]}=7'b1101011; 
        endcase
        case(seconds1)
            4'b0000: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1111101;
            4'b0001: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1100000; 
            4'b0010: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b0110111;
            4'b0011: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1100111;
            4'b0100: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1101010;
            4'b0101: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1001111;
            /*
            4'b0110: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1111100;
            4'b0111: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1000011;
            4'b1000: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1111111;
            4'b1001: {s[6],s[5],s[4],s[3],s[2],s[1],s[0]}=7'b1101011; 
            */
        endcase
        case(seconds0)
            4'b0000: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1111101;
            4'b0001: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1100000; 
            4'b0010: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b0110111;
            4'b0011: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1100111;
            4'b0100: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1101010;
            4'b0101: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1001111;
            4'b0110: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1011111;
            4'b0111: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1100001;
            4'b1000: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1111111;
            4'b1001: {s[13],s[12],s[11],s[10],s[9],s[8],s[7]}=7'b1101011; 
        endcase
        
        case(milliseconds2)
            4'b0000: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1111101;
            4'b0001: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1100000; 
            4'b0010: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b0110111;
            4'b0011: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1100111;
            4'b0100: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1101010;
            4'b0101: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1001111;
            4'b0110: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1011111;
            4'b0111: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1100001;
            4'b1000: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1111111;
            4'b1001: {k[6],k[5],k[4],k[3],k[2],k[1],k[0]}=7'b1101011;
        endcase
        case(milliseconds1)
            4'b0000: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1111101;
            4'b0001: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1100000; 
            4'b0010: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b0110111;
            4'b0011: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1100111;
            4'b0100: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1101010;
            4'b0101: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1001111;
            4'b0110: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1011111;
            4'b0111: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1100001;
            4'b1000: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1111111;
            4'b1001: {k[13],k[12],k[11],k[10],k[9],k[8],k[7]}=7'b1101011;
        endcase
        case(milliseconds0)
            4'b0000: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1111101;
            4'b0001: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1100000; 
            4'b0010: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b0110111;
            4'b0011: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1100111;
            4'b0100: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1101010;
            4'b0101: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1001111;
            4'b0110: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1011111;
            4'b0111: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1100001;
            4'b1000: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1111111;
            4'b1001: {k[20],k[19],k[18],k[17],k[16],k[15],k[14]}=7'b1101011;
        endcase
            
    end
endmodule
